`ifndef SETTINGS
`define SETTINGS

  `define COMPONENT_STRUCTURE_VERBOSITY UVM_MEDIUM
  
`endif