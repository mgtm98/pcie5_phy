`ifndef SETTINGS
`define SETTINGS

  `define COMPONENT_STRUCTURE_VERBOSITY UVM_MEDIUM
  `define PIPE_WIDTH                    32
`endif