`ifndef SETTINGS
`define SETTINGS

  `define COMPONENT_STRUCTURE_VERBOSITY UVM_MEDIUM
  `define PIPE_WIDTH                    32
  
  `define LPIF_BUS_WIDTH                512
`endif