class pipe_link_up_seq extends pipe_base_seq;

  `uvm_object_utils(pipe_link_up_seq)

  ts_s ts_sent;
  ts_s tses_sent [`NUM_OF_LANES];
  ts_s tses_received [`NUM_OF_LANES];
  int idle_data_received [`NUM_OF_LANES];

  rand gen_t           max_gen_supported;
  rand bit   [7:0]     link_number;
  rand bit   [7:0]     n_fts;
  rand int             random_start_polling;
  rand int             delay_polling;

  constraint random_start_polling_c {random_start_polling inside {0, 1, 2};}
  // Methods
  extern local task detect_state;
  extern local task polling_state;
  extern local task polling_active_state;
  extern local task polling_configuration_state;
  extern local task receiving_8_ts1;
  extern local task sending_1024_ts1;
  extern local task config_state;
  extern local task config_linkwidth_start_state_upstream;
  extern local task config_linkwidth_accept_state_upstream;
  extern local task config_lanenum_wait_state_upstream;
  extern local task config_lanenum_accept_state_upstream;
  extern local task config_complete_state_upstream;
  extern local task config_idle_state_upstream;
  extern local task config_linkwidth_start_state_downstream;
  extern local task config_linkwidth_accept_state_downstream;
  extern local task config_lanenum_wait_state_downstream;
  extern local task config_lanenum_accept_state_downstream;
  extern local task config_complete_state_downstream;
  extern local task config_idle_state_downstream;
  
  // Standard UVM Methods:
  extern function new(string name = "pipe_link_up_seq");
  extern task body;
  
endclass:pipe_link_up_seq

function pipe_link_up_seq::new(string name = "pipe_link_up_seq");
  super.new(name);
endfunction
  
task pipe_link_up_seq::body;
  super.body;
  this.randomize();

  ts_sent.n_fts            = this.n_fts;
  ts_sent.lane_number      = 0;
  ts_sent.link_number      = this.link_number;
  ts_sent.use_n_fts        = 0;
  ts_sent.use_link_number  = 0;
  ts_sent.use_lane_number  = 0;
  ts_sent.max_gen_supported = this.max_gen_supported;
  ts_sent.ts_type          = TS1;

  for (int i = 0; i < `NUM_OF_LANES; i++) begin
    tses_sent[i].n_fts            = this.n_fts;
    tses_sent[i].lane_number      = i;
    tses_sent[i].link_number      = this.link_number;
    tses_sent[i].use_n_fts        = 0;
    tses_sent[i].use_link_number  = 0;
    tses_sent[i].use_lane_number  = 0;
    tses_sent[i].max_gen_supported = this.max_gen_supported;
    tses_sent[i].ts_type          = TS1;
  end

  if (random_start_polling == 2) begin
    fork
      detect_state;
      begin
        wait(pipe_agent_config_h.start_early_polling_e.triggered)
        polling_state;
      end
    join
  end
  else begin
  detect_state;
  polling_state;
  end
  config_state;
  -> pipe_agent_config_h.link_up_finished_e;
endtask: body

task pipe_link_up_seq::detect_state;
  wait(pipe_agent_config_h.receiver_detected_e.triggered);
  `uvm_info(get_type(), "Receiver detected", UVM_MEDIUM)
endtask

task pipe_link_up_seq::polling_state;
  polling_active_state;
  polling_configuration_state;
endtask

task pipe_link_up_seq::receiving_8_ts1; //Dut sending
  int rec_8_ts1 = 0;
  //check it s okay to be in task receiving
  `uvm_info("pipe_link_up_seq", "polling state started", UVM_MEDIUM)
  wait(pipe_agent_config_h.start_polling.triggered);
  while (rec_8_ts1 < 8) begin
    wait(pipe_agent_config_h.detected_tses.triggered)
      if(pipe_agent_config_h.tses_received[0].ts_type == TS1) begin
        rec_8_ts1++;
      end
    end
endtask

//check variable option compliance or loopback in ts1?
task pipe_link_up_seq::sending_1024_ts1;
  int send_1024_ts1; 
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item");
  for (send_1024_ts1 = 0; send_1024_ts1 < 1024; send_1024_ts1++) begin
  start_item (pipe_seq_item_h);
    if (!pipe_seq_item_h.randomize() with {pipe_operation == SEND_TS; ts_sent.ts_type == TS1;})
    begin
      `uvm_error(get_name(), "Can't randomize sequence item and send TS1s")
    end
  finish_item (pipe_seq_item_h);
  end
endtask

task pipe_link_up_seq::polling_active_state;
  if (random_start_polling == 1) begin
    repeat(delay_polling) @(posedge pclk);
  end
  fork
    begin
      receiving_8_ts1;
    end
    begin
      sending_1024_ts1;
    end
  join
endtask

task pipe_link_up_seq::polling_configuration_state;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item");
  wait(pipe_agent_config_h.detected_tses.triggered)
  while (pipe_agent_config_h.tses_received[0].ts_type == TS1) begin
    start_item (pipe_seq_item_h);
        if (!pipe_seq_item_h.randomize() with {pipe_operation == SEND_TS; & ts_sent.ts_type == TS2})
        begin
          `uvm_error(get_name(), "Can't randomize sequence item and send TS1s")
        end
    finish_item (pipe_seq_item_h);
    wait(pipe_agent_config_h.detected_tses.triggered)
  end
  int rec_8_ts2 = 0;
  fork
    begin
      while(rec_8_ts2 < 8) begin
      wait(pipe_agent_config_h.detected_tses.triggered)
      if(pipe_agent_config_h.tses_received[0].ts_type == TS2) begin
        rec_8_ts2++;
      end
      end
    end
  
    begin
      for (i = 0; i < 16; i++) begin
      start_item (pipe_seq_item_h);
      if (!pipe_seq_item_h.randomize() with {pipe_operation == SEND_TS; & ts_sent.ts_type == TS2})
      begin
        `uvm_error(get_name(), "Can't randomize sequence item and send TS1s")
      end
      finish_item (pipe_seq_item_h);
      end
    end
    join
endtask

task pipe_link_up_seq::config_state;
  // Upstream
  config_linkwidth_start_state_upstream;
  config_linkwidth_accept_state_upstream;
  config_lanenum_wait_state_upstream;
  config_complete_state_upstream;
  config_idle_state_upstream;
  // Downstream
  // config_linkwidth_start_state_downstream;
  // config_linkwidth_accept_state_downstream;
  // config_lanenum_wait_state_downstream;
  // config_complete_state_downstream;
  // config_idle_state_downstream;
endtask

task pipe_link_up_seq::config_linkwidth_start_state_upstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  pipe_seq_item_h.tses_sent = tses_sent;
  int unsigned num_of_ts1s_with_non_pad_link_number [`NUM_OF_LANES];
  // Initialize the num_of_ts2_received array with zeros
  foreach(num_of_ts1s_with_non_pad_link_number[i])
  begin
    num_of_ts1s_with_non_pad_link_number[i] = 0;
  end
  // Transmit TS1s until 2 consecutive TS2s are received
  bit two_consecutive_ts1s_with_non_pad_link_number_detected = 0;
  fork
    begin
      while (!two_consecutive_ts1s_with_non_pad_link_number_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!two_consecutive_ts1s_with_non_pad_link_number_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        foreach(tses_received[i])
        begin
          if(tses_received[i].ts_type == TS1 && tses_received[i].use_link_number)
          begin
            num_of_ts1s_with_non_pad_link_number[i] += 1;
          end
          else
          begin
            num_of_ts1s_with_non_pad_link_number[i] = 0;
          end
        end
        // Check if any lane detected 2 consecutive ts2s
        foreach(num_of_ts1s_with_non_pad_link_number[i])
        begin
          if(num_of_ts1s_with_non_pad_link_number[i] == 2)
          begin
            two_consecutive_ts1s_with_non_pad_link_number_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_linkwidth_accept_state_upstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  // Use the link number of the ts1s on the first lane to be transmitted
  bit [7:0] used_link_num = tses_received[0].link_number;
  foreach(tses_sent[i])
  begin
    tses_sent[i].link_number = used_link_num;
    tses_sent[i].use_link_number = 1;
    tses_sent[i].use_lane_number = 0;
  end
  pipe_seq_item_h.tses_sent = tses_sent;
  // Send ts1s with this link number until some ts1s are received with non PAD lane number
  ts1_with_non_pad_lane_number_detected = 0;
  fork
    begin
      while (!ts1_with_non_pad_lane_number_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end
    begin
      while (!ts1_with_non_pad_lane_number_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        // Check if any ts1 received has a non PAD lane number
        foreach(tses_received[i])
        begin
          // Make sure the tses received are ts1s
          assert (tses_received[i].ts_type == TS1) 
          else   `uvm_error(get_name(), "Expected TS1s but detected TS2s")
          // Non PAD lane number
          if(tses_received[i].use_lane_num)
          begin
            ts1_with_non_pad_lane_number_detected = 1
          end
        end
      end
    end
  join
  // Get the lane numbers from the received ts1s
  foreach(tses_received[i])
  begin
    assert (tses_received[i].lane_number == i) 
    else   `uvm_error(get_name(), "the order of lane numbers are incorrect")
    tses_sent[i].lane_number = tses_received[i].lane_number;
    tses_sent[i].use_lane_number = 1;
  end
endtask

task pipe_link_up_seq::config_lanenum_wait_state_upstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  pipe_seq_item_h.tses_sent = tses_sent;
  int num_of_ts2_received [`NUM_OF_LANES];
  // Initialize the num_of_ts2_received array with zeros
  foreach(num_of_ts2_received[i])
  begin
    num_of_ts2_received[i] = 0;
  end
  // Transmit TS1s until 2 consecutive TS2s are received
  bit two_consecutive_ts2s_detected = 0;
  fork
    begin
      while (!two_consecutive_ts2s_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!two_consecutive_ts2s_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        foreach(tses_received[i])
        begin
          if(tses_received[i].ts_type == TS2)
          begin
            num_of_ts2_received[i] += 1;
          end
          else
          begin
            num_of_ts2_received[i] = 0;
          end
        end
        // Check if any lane detected 2 consecutive ts2s
        foreach(num_of_ts2_received[i])
        begin
          if(num_of_ts2_received[i] == 2)
          begin
            two_consecutive_ts2s_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_complete_state_upstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  int num_of_ts2_received [`NUM_OF_LANES];  

  // Initialize the num_of_ts2_received array with zeros
  foreach(num_of_ts2_received[i])
  begin
    num_of_ts2_received[i] = 0;
  end

  foreach (tses_sent) begin
    tses_sent.ts_type = TS2;
  end
  
  pipe_seq_item_h.tses_sent = tses_sent;

  // Transmit 16 TS2s until 8 consecutive TS2s are received
  bit eight_consecutive_ts2s_detected = 0;
  fork
    begin
      @(pipe_agent_config_h.detected_tses_e);

      for (i = 0; i < 16; i++)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end

      while (!eight_consecutive_ts2s_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!eight_consecutive_ts2s_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        
        foreach(tses_received[i])
        begin
          if(tses_received[i].ts_type == TS2)
          begin
            num_of_ts2_received[i] += 1;
          end
          else
          begin
            num_of_ts2_received[i] = 0;
          end
        end

        // Check if any lane detected 8 consecutive ts2s
        foreach(num_of_ts2_received[i])
        begin
          if(num_of_ts2_received[i] == 8)
          begin
            eight_consecutive_ts2s_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_idle_state_upstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_IDLE_DATA;
  int num_of_idle_data_received [`NUM_OF_LANES];  

  // Initialize the num_of_idle_data_received array with zeros
  foreach(num_of_idle_data_received[i])
  begin
    num_of_idle_data_received[i] = 0;
  end

  // Transmit 16 idle data until 8 consecutive idle data are received
  bit eight_consecutive_idle_data_detected = 0;
  fork
    begin
      @(pipe_agent_config_h.idle_data_detected_e);

      for (i = 0; i < 16; i++)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!eight_consecutive_idle_data_detected)
      begin
        @(pipe_agent_config_h.idle_data_detected_e);
        
        foreach(idle_data_received[i])
        begin
          begin
            num_of_idle_data_received[i] += 1;
          end
        end

        // Check if any lane detected 8 consecutive idle data
        foreach(num_of_idle_data_received[i])
        begin
          if(num_of_idle_data_received[i] == 8)
          begin
            eight_consecutive_idle_data_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_linkwidth_start_state_downstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  foreach(tses_sent[i])
  begin
    tses_sent[i].link_number = link_number;
    tses_sent[i].use_link_number = 1;
  end
  pipe_seq_item_h.tses_sent = tses_sent;
  int unsigned num_of_detected_ts1s_with_same_link_number [`NUM_OF_LANES];  
  // Initialize the num_of_detected_ts1s_with_same_link_number array with zeros
  foreach(num_of_detected_ts1s_with_same_link_number[i])
  begin
    num_of_detected_ts1s_with_same_link_number[i] = 0;
  end
  // Send ts1s with the generated link number until two ts1s are received with the same link number
  two_ts1s_with_same_link_number_detected = 0;
  fork
    begin
      while (!two_ts1s_with_same_link_number_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end
    begin
      while (!two_ts1s_with_same_link_number_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        
        foreach(tses_received[i])
        begin
          if(tses_received[i].link_number == link_number && tses_received.use_link_number)
          begin
            num_of_detected_ts1s_with_same_link_number[i] += 1;
          end
          else
          begin
            num_of_detected_ts1s_with_same_link_number[i] = 0;
          end
        end

        // Check if any lane detected 2 cosecutive ts1s with the same link number
        foreach(num_of_detected_ts1s_with_same_link_number[i])
        begin
          if(num_of_detected_ts1s_with_same_link_number[i] == 2)
          begin
            two_ts1s_with_same_link_number_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_linkwidth_accept_state_downstream;
  // Update the lane numbers to start with zero and increase sequentially
  foreach(tses_sent[i])
  begin
    tses_sent[i].lane_number = i;
    tses_sent[i].use_lane_number = 1;
  end
endtask

task pipe_link_up_seq::config_lanenum_wait_state_downstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  pipe_seq_item_h.tses_sent = tses_sent;
  int unsigned num_of_detected_ts1s_with_same_lane_numbers = 0;
  // Send ts1s with the generated lane numbers until two ts1s are received with the same link numbers
  bit two_ts1s_with_same_lane_numbers_detected = 0;
  fork
    begin
      while (!two_ts1s_with_same_lane_numbers_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end
    begin
      while (!two_ts1s_with_same_lane_numbers_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        
        bit all_lane_numbers_are_correct = 1;
        foreach(tses_received[i])
        begin
          if(tses_received[i].lane_number != tses_sent[i].lane_number || !tses_received[i].use_lane_number)
          begin
            all_lane_numbers_are_correct = 0;
          end
        end
        if (all_lane_numbers_are_correct)
        begin
          num_of_detected_ts1s_with_same_lane_numbers += 1;
        end
        else
        begin
          num_of_detected_ts1s_with_same_lane_numbers = 0;
        end

        // Check if all lane detected 2 cosecutive ts1s with the same lane numbers
        if(num_of_detected_ts1s_with_same_lane_numbers == 2)
        begin
          two_ts1s_with_same_lane_numbers_detected = 1;
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_complete_state_downstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_TSES;
  int num_of_ts2_received [`NUM_OF_LANES];  

  // Initialize the num_of_ts2_received array with zeros
  foreach(num_of_ts2_received[i])
  begin
    num_of_ts2_received[i] = 0;
  end

  foreach (tses_sent)
    tses_sent.ts_type = TS2;
  end
  
  pipe_seq_item_h.tses_sent = tses_sent;

  // Transmit 16 TS2s until 8 consecutive TS2s are received
  bit eight_consecutive_ts2s_detected = 0;
  fork
    begin
      @(pipe_agent_config_h.detected_tses_e);

      for (i = 0; i < 16; i++)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end

      while (!eight_consecutive_ts2s_detected)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!eight_consecutive_ts2s_detected)
      begin
        @(pipe_agent_config_h.detected_tses_e);
        tses_received = pipe_agent_config_h.tses_received;
        
        foreach(tses_received[i])
        begin
          if(tses_received[i].ts_type == TS2)
          begin
            num_of_ts2_received[i] += 1;
          end
          else
          begin
            num_of_ts2_received[i] = 0;
          end
        end

        // Check if any lane detected 8 consecutive ts2s
        foreach(num_of_ts2_received[i])
        begin
          if(num_of_ts2_received[i] == 8)
          begin
            eight_consecutive_ts2s_detected = 1;
          end
        end
      end
    end
  join
endtask

task pipe_link_up_seq::config_idle_state_downstream;
  pipe_seq_item pipe_seq_item_h = pipe_seq_item::type_id::create("pipe_seq_item_h");
  pipe_seq_item_h.pipe_operation = SEND_IDLE_DATA;
  int num_of_idle_data_received [`NUM_OF_LANES];  

  // Initialize the num_of_idle_data_received array with zeros
  foreach(num_of_idle_data_received[i])
  begin
    num_of_idle_data_received[i] = 0;
  end

  // Transmit 16 idle data until 8 consecutive idle data are received
  bit eight_consecutive_idle_data_detected = 0;
  fork
    begin
      @(pipe_agent_config_h.idle_data_detected_e);

      for (i = 0; i < 16; i++)
      begin
        start_item(pipe_seq_item_h);
        finish_item(pipe_seq_item_h);
      end
    end

    begin
      while (!eight_consecutive_idle_data_detected)
      begin
        @(pipe_agent_config_h.idle_data_detected_e);
        
        foreach(idle_data_received[i])
        begin
          begin
            num_of_idle_data_received[i] += 1;
          end
        end

        // Check if any lane detected 8 consecutive idle data
        foreach(num_of_idle_data_received[i])
        begin
          if(num_of_idle_data_received[i] == 8)
          begin
            eight_consecutive_idle_data_detected = 1;
          end
        end
      end
    end
  join
endtask
