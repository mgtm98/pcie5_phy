class pcie_test extends uvm_test;

  // UVM Factory Registration Macro
  //
  `uvm_component_utils(pcie_test)

  //------------------------------------------
  // Data Members
  //------------------------------------------

  //------------------------------------------
  // Component Members
  //------------------------------------------
  // The environment class
  pcie_env pcie_env_h;

  // Configuration objects

  //------------------------------------------
  // Methods
  //------------------------------------------

  // Standard UVM Methods:
  extern function new(string name = "pcie_test", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);

endclass: pcie_test

function pcie_test_test_base::new(string name = "pcie_test", uvm_component parent = null);
  super.new(name, parent);
endfunction

function void pcie_test::build_phase(uvm_phase phase);
  // env configuration
  pcie_env_config pcie_env_config_h = pcie_env_config::type_id::create("pcie_env_config_h");

  // lpif & pipe configuration creation
  lpif_agent_config lpif_agent_config_h = lpif_agent_config::type_id::create("lpif_agent_config_h");
  pipe_agent_config pipe_agent_config_h = pipe_agent_config::type_id::create("pipe_agent_config_h");

  //setting the lpif_agent conifgurations and needed handles
  if (!uvm_config_db #(virtual lpif_monitor_bfm)::get(this, "", "lpif_monitor_bfm_h", lpif_agent_config_h.lpif_monitor_bfm_h))
    `uvm_fatal("VIF CONFIG", "Cannot get() BFM interface lpif_monitor_bfm_h from uvm_config_db. Have you set() it?")
  if (!uvm_config_db #(virtual lpif_driver_bfm) ::get(this, "", "lpif_driver_bfm_h", lpif_agent_config_h.lpif_driver_bfm_h))
    `uvm_fatal("VIF CONFIG", "Cannot get() BFM interface lpif_driver_bfm_h from uvm_config_db. Have you set() it?")

  pcie_env_config_h.lpif_agent_config_h = lpif_agent_config_h;

  //setting the pipe_agent conifgurations and needed handles
  if (!uvm_config_db #(virtual pipe_monitor_bfm)::get(this, "", "pipe_monitor_bfm_h", pipe_agent_config_h.pipe_monitor_bfm_h))
    `uvm_fatal("VIF CONFIG", "Cannot get() BFM interface pipe_monitor_bfm_h from uvm_config_db. Have you set() it?")
  if (!uvm_config_db #(virtual pipe_driver_bfm) ::get(this, "", "pipe_driver_bfm_h", pipe_agent_config_h.pipe_driver_bfm_h))
    `uvm_fatal("VIF CONFIG", "Cannot get() BFM interface pipe_driver_bfm_h from uvm_config_db. Have you set() it?")

  pcie_env_config_h.pipe_agent_config_h = pipe_agent_config_h;


  
  uvm_config_db #(pcie_env_config)::set(this, "", "pcie_env_config", pcie_env_config_h);
  pcie_env_h = pcie_env::type_id::create("pcie_env_h", this);
endfunction: build_phase


task pcie_test::run_phase(uvm_phase phase);

  //get a string from the commandline arguments
  uvm_cmdline_processor cmdline_proc = uvm_cmdline_processor::get_inst();
  string arguments_value = "base_vseq"; //default value needs to be reviewed default value
  cmdline_proc.get_arg_value("+VSEQ=", arguments_value);
  string used_vsequences[$]
  uvm_split_string(arguments_value, ",", used_vsequences);

  phase.raise_objection(this, "pcie_test");

  foreach (used_vsequences[ii]) 
  begin
      //checking which vseq should be used
    case(used_vsequences[ii])
      "base_vseq":
        base_vseq vseq = base_vseq::type_id::create("vseq");
      "link_up_vseq":
        link_up_vseq vseq = link_up_vseq::type_id::create("vseq");
      "data_exchange_vseq":
        data_exchange_vseq vseq = data_exchange_vseq::type_id::create("vseq");
      "reset_vseq":
        reset_vseq vseq = reset_vseq::type_id::create("vseq");
      "enter_recovery_vseq":
        enter_recovery_vseq vseq = enter_recovery_vseq::type_id::create("vseq");
      "enter_l0s_vseq":
        enter_l0s_vseq vseq = enter_l0s_vseq::type_id::create("vseq");
      "exit_l0s_vseq":
        exit_l0s_vseq vseq = exit_l0s_vseq::type_id::create("vseq");
      "speed_change_vseq":
        speed_change_vseq vseq = speed_change_vseq::type_id::create("vseq");
    endcase

    //assigning the secquencers handles
    vseq.lpif_sequencer_h = pcie_env_h.lpif_agent_h.lpif_sequencer_h;
    vseq.pipe_sequencer_h = pcie_env_h.pipe_agent_h.pipe_sequencer_h;
    vseq.start(null); // null because no target sequencer
  end

  phase.drop_objection(this, "pcie_test");

endtask: run_phase