`ifndef SETTINGS
`define SETTINGS

  /********************** Verbosity Level Settings *************************************/
  `define COMPONENT_STRUCTURE_VERBOSITY UVM_MEDIUM
  /*************************************************************************************/
  
  /**************************** PIPE Agent Settings ************************************/
  `define PIPE_MAX_WIDTH                32
  `define PCIE_LANE_NUMBER              2
  /*************************************************************************************/

  /**************************** LPIF Agent Settings ************************************/
  `define LPIF_BUS_WIDTH                512
  /************************************************************************************/

`endif