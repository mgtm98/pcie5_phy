package utility_pkg;

	import uvm_pkg::*;
	
	`include "settings.svh"
	`include "uvm_macros.svh"
	`include "reporter.svh"
endpackage : utility_pkg