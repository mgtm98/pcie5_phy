`ifndef __PIPE_TYPES_SVH
`define __PIPE_TYPES_SVH

typedef struct 
{
  logic nothing;
} tlp_s;

typedef struct
{
  bit nothing2;
} dllp_s;

typedef enum
{
  s1
} state_e;

typedef enum
{
  s2
} speed_mode_e;

`endif


