module hvl_top;
  
  import uvm_pkg::*;
  import utility_pkg::*;
  import pcie_test_pkg::*;
  
  reporter reporter_h;
  initial begin
  	reporter_h = new();
    run_test();
  end
  
endmodule: hvl_top
  
  