package common_pkg;

  typedef bit [7:0] dllp_t [0:5];
  typedef bit [7:0] tlp_t [];

endpackage: common_pkg
