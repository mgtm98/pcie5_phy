package common_pkg;

  // TLP and DLLP definitions
  typedef bit [7:0] dllp_t [5:0];
  typedef bit [7:0] tlp_t [];

endpackage: common_pkg
