module hvl_top;
  
  import uvm_pkg::*;
  import pcie_test_pkg::*;
  
  initial begin
    run_test();
  end
  
endmodule: hvl_top
  
  