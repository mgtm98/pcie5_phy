package pcie_test_pkg;

  import uvm_pkg::*;
  import lpif_agent_pkg::*;
  import pipe_agent_pkg::*;
  import pcie_env_pkg::*;
  import pcie_seq_pkg::*;

  `include "uvm_macros.svh"  
  `include "pcie_test.svh"
  
endpackage: pcie_test_pkg
  
  